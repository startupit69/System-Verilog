import lc3b_types::*;

module cache_control
(




);

endmodule : cache_control