import lc3b_types::*;

module cache
(
	
);

cache_controller cache_controller
(

	
);

cache_datapath cache_datapath
(


);

endmodule : cache