import lc3b_types::*;
/**
 * module branch_target_adder
 * Description: computes the branch target address
 * Inputs: 
 * Outputs: br_add_out - address computed
 *
 */
 
 module br_add
(
	input lc3b_word pc_out,
	input adj9_out adj9, 
	output lc3b_word br_add_out
);

always_comb
begin

end
endmodule:br_add